module memctrl(
    input wire clk_in,  // system clock signal
    input wire rst_in,  // reset signal
    input wire rdy_in,  // ready signal, pause cpu when low

    input wire clear,

    // from to ram
    output wire

    // from ifetcher
    input wire [31:0] inst_addr,


);

endmodule